-- Steuerung