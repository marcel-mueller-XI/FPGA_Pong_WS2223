--myPack

package myPack is
type STATE_TYPE is (start, nAnB, nAnB_out, AnB_Ae, nAB_Ae, AnB_Be, nAB_Be, AB, AB_out ); 	--! mealy Automat Zustände
									--AnB_Ae bedeutet A=1 B=0 und A'event
end myPack;

package body myPack is
	
end myPack;