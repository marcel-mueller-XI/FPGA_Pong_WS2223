-- Control